`timescale  1ns/1ns
 

module  vga_pic
(
    input   wire            vga_clk     ,   //输入工作时钟,频率25MHz
    input   wire            sys_rst_n   ,   //输入复位信号,低电平有效
    input   wire    [9:0]   pix_x       ,   //输入有效显示区域像素点X轴坐标
    input   wire    [9:0]   pix_y       ,   //输入有效显示区域像素点Y轴坐标

    output  reg     [15:0]  pix_data        //输出像素点色彩信息
);

 
parameter   CHAR_B_H=   10'd192 ,   //字符开始X轴坐标
            CHAR_B_V=   10'd208 ;   //字符开始Y轴坐标

parameter   CHAR_W  =   10'd256 ,   //字符宽度
            CHAR_H  =   10'd64  ;   //字符高度

parameter   BLACK   =   16'h0000,   //黑色
            WHITE   =   16'hFFFF,   //白色
            GOLDEN  =   16'hFEC0;   //金色

//wire  define
wire    [9:0]   char_x  ;   //字符显示X轴坐标
wire    [9:0]   char_y  ;   //字符显示Y轴坐标

//reg   define
reg     [255:0] char    [31:0]  ;   //字符数据


assign  char_x  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_x - CHAR_B_H) : 10'h3FF;
assign  char_y  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_y - CHAR_B_V) : 10'h3FF;

//char:字符数据
always@(posedge vga_clk)
    begin
        char[0]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[1]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[2]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[3]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[4]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[5]     <=  256'hFC001FE07FE01FC0007F80001FFFFF801C001F000F00020001FFE2001FFFFF80;
        char[6]     <=  256'h1E001F000F0002000780FE001C0F03C01E001F000F0002000E003E00380F01C0;
        char[7]     <=  256'h1E003F000F0002000C001E00300F00C01E003F000F0002001C000F00300F00C0;
        char[8]     <=  256'h1F003F000F00020018000700200F00401F003F000F00020038000300600F0060;
        char[9]     <=  256'h1F006F000F00020038000300600F00201F006F000F00020038000100000F0000;
        char[10]    <=  256'h17006F000F00020038000000000F000017806F000F0002003C000000000F0000;
        char[11]    <=  256'h1780CF000F0002003E000000000F00001780CF000F0002001F000000000F0000;
        char[12]    <=  256'h1380CF000F0002001FC00000000F000013C0CF000F0002000FF00000000F0000;
        char[13]    <=  256'h13C18F000F00020003FE0000000F000013C18F000F00020001FF8000000F0000;
        char[14]    <=  256'h13C18F000F000200007FE000000F000011C18F000F000200001FF000000F0000;
        char[15]    <=  256'h11E30F000F0002000007FC00000F000011E30F000F0002000001FE00000F0000;
        char[16]    <=  256'h11E30F000F00020000007E00000F000010E30F000F00020000003F00000F0000;
        char[17]    <=  256'h10F30F000F00020000001F00000F000010F60F000F00020000000F80000F0000;
        char[18]    <=  256'h10F60F000F00020020000780000F000010760F000F00020030000780000F0000;
        char[19]    <=  256'h107E0F000F00020030000780000F0000107C0F000F00020010000780000F0000;
        char[20]    <=  256'h107C0F000F00020018000780000F0000103C0F000F0006001C000700000F0000;
        char[21]    <=  256'h103C0F00078004001C000F00000F000010380F0007800C001E000E00000F0000;
        char[22]    <=  256'h10380F0003C018001F001E00000F000010380F0001F070001FE07C00000F0000;
        char[23]    <=  256'h10180F0000FFE000087FF000000F0000FE107FE0003F8000001FC00000FFF000;
        char[24]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[25]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[26]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[27]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[28]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[29]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[30]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[31]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
 

    end

//pix_data:输出像素点色彩信息,根据当前像素点坐标指定当前像素点颜色数据
always@(posedge vga_clk or negedge sys_rst_n)
    if(sys_rst_n == 1'b0)
        pix_data    <= BLACK;
    else    if((((pix_x >= (CHAR_B_H - 1'b1))
                && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
                && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                && (char[char_y][10'd255 - char_x] == 1'b1))
        pix_data    <=  GOLDEN;
    else
        pix_data    <=  BLACK;

endmodule
